* Proof-of-concept circut to simulate ATmega8A microcontroller
* with N-Channel and P-Channel FETs switch.

* -----------------------------------------------------------------------------
* Including model files
* -----------------------------------------------------------------------------
.include NTA4153N.REV0.LIB
.include NTR0202PL.REV0.LIB

* -----------------------------------------------------------------------------
* Microcontroller clock (16 MHz)
* -----------------------------------------------------------------------------
Aclk_io 0 clk_io clk_iom
.model clk_iom d_osc (cntl_array=[0 1] freq_array=[16.000e6 16.000e6])

* -----------------------------------------------------------------------------
* Convert digital signals of the microcontroller to V.
* -----------------------------------------------------------------------------
Abridge [b3] [ab3] ab3_bridge
.model ab3_bridge dac_bridge (out_low=0.1 out_high=3.3)

* -----------------------------------------------------------------------------
* Microcontroller ATmega8A
* -----------------------------------------------------------------------------
.model m8a msim_m8a (config_file="pb3-pwm.conf")
Am8a clk_io -
+ [-]
+ [b0 b1 b2 b3 b4 b5 b6 b7]
+ [-] [-] [-] [-] m8a

* -----------------------------------------------------------------------------
* Switch built on n-fet and p-fet
* -----------------------------------------------------------------------------
R1	0 ab3		100k
R2	2 3		100k
R3	4 0		100k
C1	4 0		1p
XQ1	2 ab3 0		nta4153n
XQ2	4 2 3		ntr0202plt1
VDD	3 0		pwl (0 0 0ms 0 0ms 12.0v 20ms 12.0v)

* -----------------------------------------------------------------------------
* Transient analysis (step, stop, [start])
* -----------------------------------------------------------------------------
* NOTE: Step is a period which matches a frequency of 32 MHz.
.tran 31250ps 14ms

* -----------------------------------------------------------------------------
* Defining the run-time control functions
* -----------------------------------------------------------------------------
.control
run

* -----------------------------------------------------------------------------
* Plotting input and output voltages
* -----------------------------------------------------------------------------
plot v(ab3) v(4)
.endc
.end
