* PWM-to-sine converter based on ATmega8A microcontroller

* -----------------------------------------------------------------------------
* Microcontroller clock (16 MHz)
* -----------------------------------------------------------------------------
Aclk_io 0 clk_io clk_iom
.model clk_iom d_osc (cntl_array=[0 1] freq_array=[16.000e6 16.000e6])

* -----------------------------------------------------------------------------
* Microcontroller ATmega8A
* -----------------------------------------------------------------------------
.model m8a msim_m8a (config_file="firmware.conf")
Am8a clk_io -
+ [-]
+ [b0 b1 b2 b3 b4 b5 b6 b7]
+ [-] [-] [-] [-] m8a

* -----------------------------------------------------------------------------
* Convert digital signals of the microcontroller to V.
* -----------------------------------------------------------------------------
Abridge [b3] [in] ab3_bridge
.model ab3_bridge dac_bridge (out_low=0.1 out_high=3.3)

* -----------------------------------------------------------------------------
* OpAmp (to filter out all of the harmonics from a PWM signal, i.e.
*        to keep a DC component of the signal only)
* -----------------------------------------------------------------------------
.subckt opamp plus minus out
r1 plus minus 300k
a1 %vd (plus minus) outint lim
.model lim limit (out_lower_limit = -12 out_upper_limit = 12
+ fraction = true limit_range = 0.2 gain=300e3)
r3 outint out 50.0
r2 out 0 1e12
.ends opamp

* -----------------------------------------------------------------------------
* Low-pass filter (Butterworth, 3rd order, Fc = 500Hz)
*
* This filter should generally be enough to filter out all of the PWM harmonics
* starting from the ~3.9kHz carry frequency.
* -----------------------------------------------------------------------------
C2	1 0		68n
C4	2 out		100n
C6	3 0		10n
R1	in 1		5.85k
R3	1 2		9.52k
R5	2 3		8.52k
Xamp	3 out out	opamp

* -----------------------------------------------------------------------------
* Transient analysis (step, stop, [start])
* -----------------------------------------------------------------------------
* NOTE: Step is a period which matches a frequency of 32 MHz.
.tran 31250ps 14ms

* -----------------------------------------------------------------------------
* Defining the run-time control functions
* -----------------------------------------------------------------------------
.control
run

* -----------------------------------------------------------------------------
* Plotting input and output voltages
* -----------------------------------------------------------------------------
plot v(in) v(out)
.endc
.end
